// GENERATE INPLACE BEGIN head()
// GENERATE INPLACE END head



// GENERATE INPLACE BEGIN tail()
// GENERATE INPLACE END tail
